
module downsampler(
			input_data,
			output_data
			);
			
			